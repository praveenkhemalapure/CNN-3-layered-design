module table1(indx,tv);

input [4:0] indx;
output [15:0] tv;
reg [15:0] _tv;
assign tv=_tv;

always @(*) 
begin
case(indx)
0  : _tv=16'b0011001100110000;
1  : _tv=16'b0011011101100000;
2  : _tv=16'b0011100011110000;
3  : _tv=16'b0011001100110000;
4  : _tv=16'b0011011011110000;
5  : _tv=16'b0011011101100000;
6  : _tv=16'b0011100011110000;
7  : _tv=16'b0011010111000000;
8  : _tv=16'b0011011101100000;
9  : _tv=16'b0011100011110000;
10 : _tv=16'b0011001100110000;
11 : _tv=16'b0011010111000000;
12 : _tv=16'b0011100000100000;
13 : _tv=16'b0011001101110000;
14 : _tv=16'b0011010111000000;
15 : _tv=16'b0011011011110000;
16 : _tv=16'b0011100011110000;
17 : _tv=16'b0011001100110000;
18 : _tv=16'b0011010111000000;
19 : _tv=16'b0011011101100000;
20 : _tv=16'b0011100011110000;
21 : _tv=16'b0011010011010000;
22 : _tv=16'b0011011010010000;
23 : _tv=16'b0011100000100000;
24 : _tv=16'b0011100110000000;
default : _tv=16'b0000000000000000;
endcase
end 
endmodule